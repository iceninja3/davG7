module paddle(
input clk, rst, btn,
output yPos //pixel position 
);



endmodule

// in top module instantiate this module two times for two paddles