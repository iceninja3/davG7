module top(
    input clk;
    input rst;

    
);



endmodule